
* Inclusão das bibliotecas
.include	./libs/pshort.lib
.include	./libs/nshort.lib


* Declaração do subcircuito do inversor CMOS
*nome do subckt e de seus terminais
.subckt	CMOS_INVERTER   IN  OUT VDD  GND 
  
* type	drain	gate	source	bulk  model	          width  length
  MP    OUT   IN    VDD     VDD   pshort_model.0  w=3u   l=0.15u
  MN	  OUT	  IN	  GND	    GND   nshort_model.0  w=1u   l=0.15u
    
.ends

.end
 