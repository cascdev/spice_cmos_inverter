magic
tech sky130A
timestamp 1715775984
<< nwell >>
rect -94 182 71 518
<< nmos >>
rect 0 25 15 125
<< pmos >>
rect 0 200 15 500
<< ndiff >>
rect -38 105 0 125
rect -38 88 -27 105
rect -10 88 0 105
rect -38 62 0 88
rect -38 45 -27 62
rect -10 45 0 62
rect -38 25 0 45
rect 15 105 53 125
rect 15 88 25 105
rect 42 88 53 105
rect 15 62 53 88
rect 15 45 25 62
rect 42 45 53 62
rect 15 25 53 45
<< pdiff >>
rect -38 467 0 500
rect -38 450 -27 467
rect -10 450 0 467
rect -38 433 0 450
rect -38 416 -27 433
rect -10 416 0 433
rect -38 399 0 416
rect -38 382 -27 399
rect -10 382 0 399
rect -38 365 0 382
rect -38 348 -27 365
rect -10 348 0 365
rect -38 331 0 348
rect -38 314 -27 331
rect -10 314 0 331
rect -38 297 0 314
rect -38 280 -27 297
rect -10 280 0 297
rect -38 263 0 280
rect -38 246 -27 263
rect -10 246 0 263
rect -38 229 0 246
rect -38 212 -27 229
rect -10 212 0 229
rect -38 200 0 212
rect 15 467 53 500
rect 15 450 25 467
rect 42 450 53 467
rect 15 433 53 450
rect 15 416 25 433
rect 42 416 53 433
rect 15 399 53 416
rect 15 382 25 399
rect 42 382 53 399
rect 15 365 53 382
rect 15 348 25 365
rect 42 348 53 365
rect 15 331 53 348
rect 15 314 25 331
rect 42 314 53 331
rect 15 297 53 314
rect 15 280 25 297
rect 42 280 53 297
rect 15 263 53 280
rect 15 246 25 263
rect 42 246 53 263
rect 15 229 53 246
rect 15 212 25 229
rect 42 212 53 229
rect 15 200 53 212
<< ndiffc >>
rect -27 88 -10 105
rect -27 45 -10 62
rect 25 88 42 105
rect 25 45 42 62
<< pdiffc >>
rect -27 450 -10 467
rect -27 416 -10 433
rect -27 382 -10 399
rect -27 348 -10 365
rect -27 314 -10 331
rect -27 280 -10 297
rect -27 246 -10 263
rect -27 212 -10 229
rect 25 450 42 467
rect 25 416 42 433
rect 25 382 42 399
rect 25 348 42 365
rect 25 314 42 331
rect 25 280 42 297
rect 25 246 42 263
rect 25 212 42 229
<< psubdiff >>
rect -76 105 -38 125
rect -76 88 -61 105
rect -44 88 -38 105
rect -76 62 -38 88
rect -76 45 -61 62
rect -44 45 -38 62
rect -76 25 -38 45
<< nsubdiff >>
rect -76 467 -38 500
rect -76 450 -61 467
rect -44 450 -38 467
rect -76 433 -38 450
rect -76 416 -61 433
rect -44 416 -38 433
rect -76 399 -38 416
rect -76 382 -61 399
rect -44 382 -38 399
rect -76 365 -38 382
rect -76 348 -61 365
rect -44 348 -38 365
rect -76 331 -38 348
rect -76 314 -61 331
rect -44 314 -38 331
rect -76 297 -38 314
rect -76 280 -61 297
rect -44 280 -38 297
rect -76 263 -38 280
rect -76 246 -61 263
rect -44 246 -38 263
rect -76 229 -38 246
rect -76 212 -61 229
rect -44 212 -38 229
rect -76 200 -38 212
<< psubdiffcont >>
rect -61 88 -44 105
rect -61 45 -44 62
<< nsubdiffcont >>
rect -61 450 -44 467
rect -61 416 -44 433
rect -61 382 -44 399
rect -61 348 -44 365
rect -61 314 -44 331
rect -61 280 -44 297
rect -61 246 -44 263
rect -61 212 -44 229
<< poly >>
rect 0 500 15 525
rect -94 168 -59 177
rect 0 168 15 200
rect -94 151 -85 168
rect -68 151 15 168
rect -94 142 -59 151
rect 0 125 15 151
rect 0 0 15 25
<< polycont >>
rect -85 151 -68 168
<< locali >>
rect -95 562 71 563
rect -78 545 -61 562
rect -44 545 -27 562
rect -10 545 7 562
rect 24 545 41 562
rect 58 545 71 562
rect -95 543 71 545
rect -61 500 -38 543
rect -61 467 -10 500
rect -44 450 -27 467
rect -61 433 -10 450
rect -44 416 -27 433
rect -61 399 -10 416
rect -44 382 -27 399
rect -61 365 -10 382
rect -44 348 -27 365
rect -61 331 -10 348
rect -44 314 -27 331
rect -61 297 -10 314
rect -44 280 -27 297
rect -61 263 -10 280
rect -44 246 -27 263
rect -61 229 -10 246
rect -44 212 -27 229
rect -61 200 -10 212
rect 25 467 42 500
rect 25 433 42 450
rect 25 399 42 416
rect 25 365 42 382
rect 25 331 42 348
rect 25 297 42 314
rect 25 263 42 280
rect 25 229 42 246
rect -94 168 -59 177
rect -94 151 -85 168
rect -68 151 -59 168
rect -94 142 -59 151
rect 25 170 42 212
rect 25 169 67 170
rect 25 152 40 169
rect 57 152 67 169
rect 25 150 67 152
rect -61 105 -10 125
rect -44 88 -27 105
rect -61 62 -10 88
rect -44 45 -27 62
rect -61 25 -10 45
rect 25 105 42 150
rect 25 62 42 88
rect 25 25 42 45
rect -61 -21 -38 25
rect -96 -22 70 -21
rect -79 -39 -61 -22
rect -44 -23 70 -22
rect -44 -39 -25 -23
rect -96 -40 -25 -39
rect -8 -40 10 -23
rect 27 -40 44 -23
rect 61 -40 70 -23
rect -96 -41 70 -40
<< viali >>
rect -95 545 -78 562
rect -61 545 -44 562
rect -27 545 -10 562
rect 7 545 24 562
rect 41 545 58 562
rect 40 152 57 169
rect -96 -39 -79 -22
rect -61 -39 -44 -22
rect -25 -40 -8 -23
rect 10 -40 27 -23
rect 44 -40 61 -23
<< metal1 >>
rect -100 562 77 568
rect -100 545 -95 562
rect -78 545 -61 562
rect -44 545 -27 562
rect -10 545 7 562
rect 24 545 41 562
rect 58 545 77 562
rect -100 538 77 545
rect 25 169 70 175
rect 25 152 40 169
rect 57 152 70 169
rect 25 145 70 152
rect -102 -22 75 -15
rect -102 -39 -96 -22
rect -79 -39 -61 -22
rect -44 -23 75 -22
rect -44 -39 -25 -23
rect -102 -40 -25 -39
rect -8 -40 10 -23
rect 27 -40 44 -23
rect 61 -40 75 -23
rect -102 -45 75 -40
<< labels >>
rlabel viali -27 545 -10 562 1 VDD
rlabel viali -25 -40 -8 -23 1 GND
rlabel polycont -85 151 -68 168 1 IN
rlabel viali 40 152 57 169 1 OUT
rlabel metal1 -102 -20 -90 -15 1 GND
rlabel metal1 55 145 67 150 1 OUT
rlabel metal1 -60 563 -48 568 5 VDD
rlabel locali -94 142 -85 177 1 IN
rlabel polycont -80 156 -74 164 1 IN
<< end >>
