* SPICE3 file created from layout_inverter.ext - technology: sky130A

* incluir libs
.include	../libs/pshort.lib
.include	../libs/nshort.lib

.subckt	cmos_inv OUT IN	VDD	GND
* type	drain	gate	source	bulk  model	           width    length
 M1000  OUT     IN      VDD     VDD   pshort_model.0   w=3e+06u l=150000u
+  ad=1.14e+12p pd=6.76e+06u as=1.14e+12p ps=6.76e+06u

M1001   OUT     IN      GND     GND   nshort_model.0   w=1e+06u l=150000u
+  ad=3.8e+11p pd=2.76e+06u as=3.8e+11p ps=2.76e+06u

.ends

.end

